// ВНИМАНИЕ!
// Можно изменять ТОЛЬКО части кода, помеченные "(*)",
//   и ТОЛЬКО так, как написано у "(*)".
module main(x, on, start, y, s, b, regime, active, clk, rst);
  // // (*) По необходимости можно добавть "reg" в объявлениях выходных точек, задающихся в управляющем автомате.
  input [7:0] x;
  input [1:0] on;
  input start;
  output [7:0] y;
  output [2:0] s;
  output b, active;
  output [1:0] regime;
  input clk, rst;
  
  // (*) По необходимости можно заменить wire на reg для любых точек далее.
  wire [1:0] y_select_next, s_step;
  wire y_en, s_en, y_upd, s_sub, s_zero;
  
  // Основная часть операционного автомата.
  datapath _datapath(
    .x(x),
    .y(y),
    .s(s),
    .b(b),
    .s_en(s_en),
    .s_step(s_step),
    .s_sub(s_sub),
    .s_zero(s_zero),
    .y_en(y_en),
    .y_select_next(y_select_next),
    .y_upd(y_upd),
    .clk(clk),
    .rst(rst)
  );
  
  // Распознавание свойств данных в операционном автомате.
  // (*) Здесь следует по необходимости объявить новые управляющие точки
  //   и реализовать задающие их подсхемы
  //   (преобразующие данные в управление).
  
  // Управляющий автомат.
  // (*) Здесь следует написать схему, основная часть которой - это
  //   типовая реализация управляющего символьного автомата,
  //   заставляющая схему main выполняться согласно условию.
endmodule
